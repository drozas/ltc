package constantes is
	constant n: natural:= 16;
end constantes;