package constantes is
	constant n: natural:= 8;
end constantes;